-- This Source Code Form is subject to the terms of the Mozilla Public
-- License, v. 2.0. If a copy of the MPL was not distributed with this file,
-- You can obtain one at http://mozilla.org/MPL/2.0/.
--
-- Copyright (c) 2014, Lars Asplund lars.anders.asplund@gmail.com

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

library vunit_lib;
context vunit_lib.vunit_context;
use vunit_lib.array_pkg.all;

entity tb_sobel_x is
  generic (
    runner_cfg : runner_cfg_t;
    data_width : natural := 14;
    output_path : string);
end entity;

architecture tb of tb_sobel_x is
  signal clk : std_logic := '0';
  signal input_tvalid : std_logic := '0';
  signal input_tlast : std_logic := '0';
  signal input_tdata : unsigned(data_width-1 downto 0) := (others => '0');
  signal output_tvalid : std_logic;
  signal output_tlast : std_logic;
  signal output_tdata : signed(input_tdata'length downto 0);

  shared variable image : array_t;
  shared variable reference_image : array_t;
  signal start, data_check_done, stimuli_done : boolean := false;
begin

  main : process
    procedure sobel_x(variable image : inout array_t;
                      variable result : inout array_t) is
    begin
      result.init_2d(width => image.width,
                     height => image.height,
                     bit_width => image.bit_width+1,
                     is_signed => true);

      for y in 0 to image.height-1 loop
        for x in 0 to image.width-1 loop
          result.set(x, y,
                     value => (image.get(minimum(x+1, image.width-1),y) -
                               image.get(maximum(x-1, 0), y)));
        end loop;
      end loop;

    end procedure;

    variable seed1 : positive := 12315;
    variable seed2 : positive := 8918239;

    procedure randomize(variable arr : inout array_t) is
      impure function random_value return integer is
        variable random_real : real;
      begin
        uniform(seed1, seed2, random_real);
        if arr.is_signed then
          random_real := random_real - 0.5;
        end if;
        return integer(trunc(random_real * 2.0**arr.bit_width));
      end function;
    begin
      for idx in 0 to arr.length-1 loop
        arr.set(idx, value => random_value);
      end loop;
    end procedure;

    procedure test_one_image(width, height : natural) is
    begin
      image.init_2d(width => width, height => height,
                    bit_width => input_tdata'length,
                    is_signed => false);
      randomize(image);
      sobel_x(image, result => reference_image);

      wait until rising_edge(clk);
      start <= true;
      wait until rising_edge(clk);
      start <= false;

      wait until (stimuli_done and
                  data_check_done and
                  rising_edge(clk));
    end procedure;

  begin
    test_runner_setup(runner, runner_cfg);
    test_one_image(128, 64);
    test_one_image(1, 13);
    test_one_image(16, 1);
    test_one_image(1, 1);
    test_runner_cleanup(runner);
    wait;
  end process;

  stimuli_process : process
  begin
    wait until start and rising_edge(clk);
    stimuli_done <= false;

    report ("Sending image of size " &
            to_string(image.width) & "x" &
            to_string(image.height));

    for y in 0 to image.height-1 loop
      for x in 0 to image.width-1 loop
        wait until rising_edge(clk);
        input_tvalid <= '1';
        input_tlast <= '1' when x = image.width-1 else '0';
        input_tdata <= to_unsigned(image.get(x,y), input_tdata'length);
      end loop;
    end loop;

    wait until rising_edge(clk);
    input_tvalid <= '0';

    stimuli_done <= true;
  end process;

  data_check_process : process
  begin
    wait until start and rising_edge(clk);
    data_check_done <= false;
    for y in 0 to reference_image.height-1 loop
      for x in 0 to reference_image.width-1 loop
        wait until output_tvalid = '1' and rising_edge(clk);
        check_equal(output_tlast, x = reference_image.width-1);
        check_equal(output_tdata, reference_image.get(x, y),
                    "x=" & to_string(x) & " y=" & to_string(y));
      end loop;
    end loop;
    report ("Done checking image of size " &
            to_string(reference_image.width) & "x" &
            to_string(reference_image.height));
    data_check_done <= true;
  end process;

  clk <= not clk after 1 ns;

  dut : entity work.sobel_x
    generic map (
      data_width => input_tdata'length)
    port map (
      clk           => clk,
      input_tvalid  => input_tvalid,
      input_tlast   => input_tlast,
      input_tdata   => input_tdata,
      output_tvalid => output_tvalid,
      output_tlast  => output_tlast,
      output_tdata  => output_tdata);

end architecture;
